-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: framebuffer.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity framebuffer is
port (
data : in std_logic_vector(15 downto 0);
wraddress : in std_logic_vector(12 downto 0);
wrclock : in std_logic;
wren : in std_logic;
rdaddress : in std_logic_vector(12 downto 0);
rdclock : in std_logic;
q : out std_logic_vector(15 downto 0)
);
end entity;

architecture rtl of framebuffer is
type ram_type is array(0 to 8191) of std_logic_vector(15 downto 0);
signal ram : ram_type := (others => (others => '0'));
signal rd_data : std_logic_vector(15 downto 0);
begin


process(wrclock)
begin
    if rising_edge(wrclock) then
        if wren = '1' then
            ram(to_integer(unsigned(wraddress))) <= data;
        end if;
    end if;
end process;


process(rdclock)
begin
    if rising_edge(rdclock) then
        rd_data <= ram(to_integer(unsigned(rdaddress)));
    end if;
end process;

q <= rd_data;

end architecture;
